-- Copyright (C) 2016  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel MegaCore Function License Agreement, or other 
-- applicable license agreement, including, without limitation, 
-- that your use is for the sole purpose of programming logic 
-- devices manufactured by Intel and sold by Intel or its 
-- authorized distributors.  Please refer to the applicable 
-- agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 16.1.0 Build 196 10/24/2016 SJ Standard Edition"
-- CREATED		"Wed Nov 01 11:46:10 2017"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY projectA IS 
	PORT
	(
		reset :  IN  STD_LOGIC;
		clock :  IN  STD_LOGIC;
		four :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END projectA;

ARCHITECTURE bdf_type OF projectA IS 

COMPONENT alu
	PORT(ALU_OP : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 i_A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 i_B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 shamt : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 zero : OUT STD_LOGIC;
		 ALU_out : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT dmem
GENERIC (depth_exp_of_2 : INTEGER;
			mif_filename : STRING
			);
	PORT(clock : IN STD_LOGIC;
		 wren : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 byteena : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT imem
GENERIC (depth_exp_of_2 : INTEGER;
			mif_filename : STRING
			);
	PORT(clock : IN STD_LOGIC;
		 wren : IN STD_LOGIC;
		 address : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
		 byteena : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 q : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT concatonate
	PORT(highFourBits : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 low28Bits : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
		 concatonated : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux21_32bit
	PORT(i_sel : IN STD_LOGIC;
		 i_0 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 i_1 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_mux : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT mux21_5bit
	PORT(i_sel : IN STD_LOGIC;
		 i_0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 i_1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 o_mux : OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
	);
END COMPONENT;

COMPONENT sll_2
	PORT(i_to_shift : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_shifted : OUT STD_LOGIC_VECTOR(27 DOWNTO 0)
	);
END COMPONENT;

COMPONENT sign_extender_16_32
	PORT(i_to_extend : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 o_extended : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT adder_32
	PORT(i_A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 i_B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_F : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT main_control
	PORT(i_instruction : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_reg_dest : OUT STD_LOGIC;
		 o_jump : OUT STD_LOGIC;
		 o_branch : OUT STD_LOGIC;
		 o_mem_to_reg : OUT STD_LOGIC;
		 o_mem_write : OUT STD_LOGIC;
		 o_ALU_src : OUT STD_LOGIC;
		 o_reg_write : OUT STD_LOGIC;
		 o_ALU_op : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

COMPONENT pc_reg
	PORT(CLK : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 i_next_PC : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 o_PC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

COMPONENT register_file
	PORT(CLK : IN STD_LOGIC;
		 w_en : IN STD_LOGIC;
		 reset : IN STD_LOGIC;
		 rs_sel : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 rt_sel : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 w_data : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		 w_sel : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		 rs_data : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		 rt_data : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	ALU_out :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	o_F :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	o_PC :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	q :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(0 TO 4);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC_VECTOR(0 TO 3);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(0 TO 31);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(27 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC_VECTOR(4 DOWNTO 0);


BEGIN 
SYNTHESIZED_WIRE_0 <= "0000";
SYNTHESIZED_WIRE_2 <= "00000";
SYNTHESIZED_WIRE_4 <= "1111";
SYNTHESIZED_WIRE_6 <= '0';
SYNTHESIZED_WIRE_7 <= "1111";
SYNTHESIZED_WIRE_8 <= "00000000000000000000000000000000";



b2v_ALU2 : alu
PORT MAP(ALU_OP => SYNTHESIZED_WIRE_0,
		 i_A => o_F,
		 i_B => SYNTHESIZED_WIRE_1,
		 shamt => SYNTHESIZED_WIRE_2,
		 ALU_out => SYNTHESIZED_WIRE_19);


b2v_dmemory : dmem
GENERIC MAP(depth_exp_of_2 => 10,
			mif_filename => "dmem.mif"
			)
PORT MAP(clock => clock,
		 wren => SYNTHESIZED_WIRE_3,
		 address => ALU_out(11 DOWNTO 2),
		 byteena => SYNTHESIZED_WIRE_4,
		 data => SYNTHESIZED_WIRE_31,
		 q => SYNTHESIZED_WIRE_25);




b2v_imemory : imem
GENERIC MAP(depth_exp_of_2 => 10,
			mif_filename => "imem.mif"
			)
PORT MAP(clock => clock,
		 wren => SYNTHESIZED_WIRE_6,
		 address => o_PC(11 DOWNTO 2),
		 byteena => SYNTHESIZED_WIRE_7,
		 data => SYNTHESIZED_WIRE_8,
		 q => q);


b2v_inst : concatonate
PORT MAP(highFourBits => o_F,
		 low28Bits => SYNTHESIZED_WIRE_9,
		 concatonated => SYNTHESIZED_WIRE_15);


b2v_inst1 : alu
PORT MAP(ALU_OP => SYNTHESIZED_WIRE_10,
		 i_A => SYNTHESIZED_WIRE_11,
		 i_B => SYNTHESIZED_WIRE_12,
		 shamt => q(10 DOWNTO 6),
		 zero => SYNTHESIZED_WIRE_17,
		 ALU_out => ALU_out);


b2v_inst11 : mux21_32bit
PORT MAP(i_sel => SYNTHESIZED_WIRE_13,
		 i_0 => SYNTHESIZED_WIRE_14,
		 i_1 => SYNTHESIZED_WIRE_15,
		 o_mux => SYNTHESIZED_WIRE_27);


SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_16 AND SYNTHESIZED_WIRE_17;



b2v_inst14 : mux21_32bit
PORT MAP(i_sel => SYNTHESIZED_WIRE_18,
		 i_0 => o_F,
		 i_1 => SYNTHESIZED_WIRE_19,
		 o_mux => SYNTHESIZED_WIRE_14);


b2v_inst17 : mux21_32bit
PORT MAP(i_sel => SYNTHESIZED_WIRE_20,
		 i_0 => SYNTHESIZED_WIRE_31,
		 i_1 => SYNTHESIZED_WIRE_32,
		 o_mux => SYNTHESIZED_WIRE_12);


b2v_inst18 : mux21_5bit
PORT MAP(i_sel => SYNTHESIZED_WIRE_23,
		 i_0 => q(20 DOWNTO 16),
		 i_1 => q(15 DOWNTO 11),
		 o_mux => SYNTHESIZED_WIRE_30);


b2v_inst2 : sll_2
PORT MAP(i_to_shift => q,
		 o_shifted => SYNTHESIZED_WIRE_9);


b2v_inst21 : mux21_32bit
PORT MAP(i_sel => SYNTHESIZED_WIRE_24,
		 i_0 => ALU_out,
		 i_1 => SYNTHESIZED_WIRE_25,
		 o_mux => SYNTHESIZED_WIRE_29);


b2v_inst22 : sign_extender_16_32
PORT MAP(i_to_extend => q(15 DOWNTO 0),
		 o_extended => SYNTHESIZED_WIRE_32);




b2v_inst3 : sll_2
PORT MAP(i_to_shift => SYNTHESIZED_WIRE_32,
		 o_shifted => SYNTHESIZED_WIRE_1);



b2v_inst999 : adder_32
PORT MAP(i_A => q,
		 i_B => four,
		 o_F => o_F);


b2v_mainControl : main_control
PORT MAP(i_instruction => q,
		 o_reg_dest => SYNTHESIZED_WIRE_23,
		 o_jump => SYNTHESIZED_WIRE_13,
		 o_branch => SYNTHESIZED_WIRE_16,
		 o_mem_to_reg => SYNTHESIZED_WIRE_24,
		 o_mem_write => SYNTHESIZED_WIRE_3,
		 o_ALU_src => SYNTHESIZED_WIRE_20,
		 o_reg_write => SYNTHESIZED_WIRE_28,
		 o_ALU_op => SYNTHESIZED_WIRE_10);


b2v_pcRegister : pc_reg
PORT MAP(CLK => clock,
		 reset => reset,
		 i_next_PC => SYNTHESIZED_WIRE_27,
		 o_PC => o_PC);


b2v_registerFile : register_file
PORT MAP(CLK => clock,
		 w_en => SYNTHESIZED_WIRE_28,
		 reset => reset,
		 rs_sel => q(15 DOWNTO 11),
		 rt_sel => q(20 DOWNTO 16),
		 w_data => SYNTHESIZED_WIRE_29,
		 w_sel => SYNTHESIZED_WIRE_30,
		 rs_data => SYNTHESIZED_WIRE_11,
		 rt_data => SYNTHESIZED_WIRE_31);


END bdf_type;